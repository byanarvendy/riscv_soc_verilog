`include "logical/rtl/core/riscv_32i.v"
`include "logical/rtl/core/register_file.v"
`include "logical/rtl/core/alu/alu.v"
`include "logical/rtl/core/alu/instruction_mux.v"
`include "logical/rtl/core/alu/rv32i/instruction_r.v"
`include "logical/rtl/core/alu/rv32i/instruction_i.v"
`include "logical/rtl/core/alu/rv32i/instruction_s.v"
`include "logical/rtl/core/alu/rv32i/instruction_b.v"
`include "logical/rtl/core/alu/rv32i/instruction_u.v"
`include "logical/rtl/core/alu/rv32i/instruction_j.v"
`include "logical/rtl/soc/ram/memory_ram.v"
`include "logical/rtl/soc/rom/memory_rom.v"
`include "logical/rtl/soc/axi4_lite/axi4_lite_master.v"
`include "logical/rtl/soc/axi4_lite/axi4_lite_slave.v"
`include "logical/rtl/soc/axi4_lite/axi4_lite_interconnect_m1s2.v"
`include "logical/rtl/soc/axi4_lite/wrapper/axi4_lite_cpu_wrapper.v"
`include "logical/rtl/soc/axi4_lite/wrapper/axi4_lite_ram_wrapper.v"
`include "logical/rtl/soc/axi4_lite/wrapper/axi4_lite_rom_wrapper.v"
`include "logical/rtl/soc/gpio/gpio.v"
`include "logical/rtl/soc/axi4_lite/wrapper/axi4_lite_gpio_wrapper.v"